interface wrapperif (
    clk
);
  input clk;
  logic MOSI, SS_n, rst_n;
  logic MISO,MISO_exp; 
endinterface
